library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

package func_pkg is
    function log2ceil(val : natural) return natural;
end func_pkg;
